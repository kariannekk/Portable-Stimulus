//====================================================================
// Created       : Karianne Krokan Kragseth at 2018-03-07
//====================================================================

package paTest_par;
  
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "par_uvm/par_sequencer.sv"
  `include "par_uvm/par_driver.sv"
  `include "par_uvm/par_monitor.sv"
  `include "par_uvm/par_agent.sv"
  `include "par_uvm/par_env.sv"

endpackage : paTest_par